//


virtual class transactor
